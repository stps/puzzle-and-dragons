import lc3b_types::*;

module dep_check_logic
(
	input logic sr1_needed,
	input logic sr2_needed,
	input lc3b_opcode opcode,
	
	input logic ex_ld_cc,
	input logic mem_ld_cc,
	input logic wb_load_cc
	
);
         always_comb
         begin
				
				
         end
endmodule : mem_stall_logic