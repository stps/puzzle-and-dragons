module execute
begin

endmodule : execute
