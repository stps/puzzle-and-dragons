module write_back
begin

endmodule : write_back
