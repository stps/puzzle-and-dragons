import lc3b_types::*;

module forwarding_unit
(
    input lc3bword ex_mem_regdata,
    input lc3bword mem_wb_regdata,
    
);