import lc3b_types::*;

module fetch
(
	input clk,
	input pc_mux_sel,

	output new_pc,
	output ir,
	output valid,
	output stall
);

endmodule : fetch